module _32_bits_and(Res, A, B);
input [31:0] A, B;
output [31:0] Res;

and A0(Res[0], A[0], B[0]);
and A1(Res[1], A[1], B[1]);
and A2(Res[2], A[2], B[2]);
and A3(Res[3], A[3], B[3]);
and A4(Res[4], A[4], B[4]);
and A5(Res[5], A[5], B[5]);
and A6(Res[6], A[6], B[6]);
and A7(Res[7], A[7], B[7]);
and A8(Res[8], A[8], B[8]);
and A9(Res[9], A[9], B[9]);
and A10(Res[10], A[10], B[10]);
and A11(Res[11], A[11], B[11]);
and A12(Res[12], A[12], B[12]);
and A13(Res[13], A[13], B[13]);
and A14(Res[14], A[14], B[14]);
and A15(Res[15], A[15], B[15]);
and A16(Res[16], A[16], B[16]);
and A17(Res[17], A[17], B[17]);
and A18(Res[18], A[18], B[18]);
and A19(Res[19], A[19], B[19]);
and A20(Res[20], A[20], B[20]);
and A21(Res[21], A[21], B[21]);
and A22(Res[22], A[22], B[22]);
and A23(Res[23], A[23], B[23]);
and A24(Res[24], A[24], B[24]);
and A25(Res[25], A[25], B[25]);
and A26(Res[26], A[26], B[26]);
and A27(Res[27], A[27], B[27]);
and A28(Res[28], A[28], B[28]);
and A29(Res[29], A[29], B[29]);
and A30(Res[30], A[30], B[30]);
and A31(Res[31], A[31], B[31]);

endmodule